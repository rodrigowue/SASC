.SUBCKT NANDD0BWP A B OUT VDD VSS
*.pininfo A:I B:I OUT:O VSS:G VDD:P
MP0 VDD A OUT VDD PCH W=5e-06 NF=1 L=4e-08
MP1 VDD B OUT VDD PCH W=5e-06 NF=1 L=4e-08
MN0 OUT A rand0 VSS NCH W=5e-06 NF=1 L=4e-08
MN1 rand0 B VSS VSS NCH W=5e-06 NF=1 L=4e-08

.ENDS

